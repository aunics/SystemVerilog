class Singleton_ex;

endclass
