class Constraint_Ex;

endclass // Constraint_Ex

module test;

initial begin
end
   
endmodule // test
