class constraint_layering;
endclass // constraint_layering

module test;

initial begin
end

endmodule // test

     
